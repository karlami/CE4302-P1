module FixedAdd #(parameter DATA_WIDTH = 16)(
    input logic [DATA_WIDTH-1:0] operand1,
    input logic [DATA_WIDTH-1:0] operand2,
    output logic [DATA_WIDTH-1:0] result
);

endmodule

